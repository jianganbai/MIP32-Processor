module InstructionMemory(reset, Address, Instruction);
	input reset;
	input [31:0] Address;
	output reg [31:0] Instruction;
	
	always @(*)
	   if(reset)
	       Instruction <= 32'h00000000;
	   else
	       case (Address[11:2])   //���2λΪ00������֧��1024�����
                10'd0: Instruction <= 32'h08000003;
           10'd1: Instruction <= 32'h08000158;
           10'd2: Instruction <= 32'h0800018b;
           10'd3: Instruction <= 32'h201f0014;
           10'd4: Instruction <= 32'h03e00008;
           10'd5: Instruction <= 32'h0000f820;
           10'd6: Instruction <= 32'h20080000;
           10'd7: Instruction <= 32'h3c094000;
           10'd8: Instruction <= 32'h21290008;
           10'd9: Instruction <= 32'had280000;
           10'd10: Instruction <= 32'h200802e2;
           10'd11: Instruction <= 32'hac080000;
           10'd12: Instruction <= 32'h2008177c;
           10'd13: Instruction <= 32'hac080004;
           10'd14: Instruction <= 32'h2008756a;
           10'd15: Instruction <= 32'hac080008;
           10'd16: Instruction <= 32'h20087d9d;
           10'd17: Instruction <= 32'hac08000c;
           10'd18: Instruction <= 32'h20085f7d;
           10'd19: Instruction <= 32'hac080010;
           10'd20: Instruction <= 32'h20086924;
           10'd21: Instruction <= 32'hac080014;
           10'd22: Instruction <= 32'h20082246;
           10'd23: Instruction <= 32'hac080018;
           10'd24: Instruction <= 32'h200808cb;
           10'd25: Instruction <= 32'hac08001c;
           10'd26: Instruction <= 32'h200822ef;
           10'd27: Instruction <= 32'hac080020;
           10'd28: Instruction <= 32'h2008211e;
           10'd29: Instruction <= 32'hac080024;
           10'd30: Instruction <= 32'h20085fb0;
           10'd31: Instruction <= 32'hac080028;
           10'd32: Instruction <= 32'h20085bcb;
           10'd33: Instruction <= 32'hac08002c;
           10'd34: Instruction <= 32'h20085673;
           10'd35: Instruction <= 32'hac080030;
           10'd36: Instruction <= 32'h20081646;
           10'd37: Instruction <= 32'hac080034;
           10'd38: Instruction <= 32'h2008115f;
           10'd39: Instruction <= 32'hac080038;
           10'd40: Instruction <= 32'h2008528a;
           10'd41: Instruction <= 32'hac08003c;
           10'd42: Instruction <= 32'h20081113;
           10'd43: Instruction <= 32'hac080040;
           10'd44: Instruction <= 32'h2008430c;
           10'd45: Instruction <= 32'hac080044;
           10'd46: Instruction <= 32'h20084953;
           10'd47: Instruction <= 32'hac080048;
           10'd48: Instruction <= 32'h20087318;
           10'd49: Instruction <= 32'hac08004c;
           10'd50: Instruction <= 32'h20084c6e;
           10'd51: Instruction <= 32'hac080050;
           10'd52: Instruction <= 32'h20085728;
           10'd53: Instruction <= 32'hac080054;
           10'd54: Instruction <= 32'h200862b7;
           10'd55: Instruction <= 32'hac080058;
           10'd56: Instruction <= 32'h20082cff;
           10'd57: Instruction <= 32'hac08005c;
           10'd58: Instruction <= 32'h200876b9;
           10'd59: Instruction <= 32'hac080060;
           10'd60: Instruction <= 32'h2008118a;
           10'd61: Instruction <= 32'hac080064;
           10'd62: Instruction <= 32'h2008440c;
           10'd63: Instruction <= 32'hac080068;
           10'd64: Instruction <= 32'h200822d4;
           10'd65: Instruction <= 32'hac08006c;
           10'd66: Instruction <= 32'h20086604;
           10'd67: Instruction <= 32'hac080070;
           10'd68: Instruction <= 32'h20087690;
           10'd69: Instruction <= 32'hac080074;
           10'd70: Instruction <= 32'h20080c84;
           10'd71: Instruction <= 32'hac080078;
           10'd72: Instruction <= 32'h2008320b;
           10'd73: Instruction <= 32'hac08007c;
           10'd74: Instruction <= 32'h200810be;
           10'd75: Instruction <= 32'hac080080;
           10'd76: Instruction <= 32'h2008367c;
           10'd77: Instruction <= 32'hac080084;
           10'd78: Instruction <= 32'h200830ac;
           10'd79: Instruction <= 32'hac080088;
           10'd80: Instruction <= 32'h20082d0f;
           10'd81: Instruction <= 32'hac08008c;
           10'd82: Instruction <= 32'h20082f7c;
           10'd83: Instruction <= 32'hac080090;
           10'd84: Instruction <= 32'h20085825;
           10'd85: Instruction <= 32'hac080094;
           10'd86: Instruction <= 32'h20084a4e;
           10'd87: Instruction <= 32'hac080098;
           10'd88: Instruction <= 32'h20087b93;
           10'd89: Instruction <= 32'hac08009c;
           10'd90: Instruction <= 32'h20082bf6;
           10'd91: Instruction <= 32'hac0800a0;
           10'd92: Instruction <= 32'h20087bed;
           10'd93: Instruction <= 32'hac0800a4;
           10'd94: Instruction <= 32'h20081f96;
           10'd95: Instruction <= 32'hac0800a8;
           10'd96: Instruction <= 32'h20081522;
           10'd97: Instruction <= 32'hac0800ac;
           10'd98: Instruction <= 32'h20080152;
           10'd99: Instruction <= 32'hac0800b0;
           10'd100: Instruction <= 32'h20084af2;
           10'd101: Instruction <= 32'hac0800b4;
           10'd102: Instruction <= 32'h20082573;
           10'd103: Instruction <= 32'hac0800b8;
           10'd104: Instruction <= 32'h200809fe;
           10'd105: Instruction <= 32'hac0800bc;
           10'd106: Instruction <= 32'h200871a6;
           10'd107: Instruction <= 32'hac0800c0;
           10'd108: Instruction <= 32'h20086689;
           10'd109: Instruction <= 32'hac0800c4;
           10'd110: Instruction <= 32'h20080140;
           10'd111: Instruction <= 32'hac0800c8;
           10'd112: Instruction <= 32'h20080e27;
           10'd113: Instruction <= 32'hac0800cc;
           10'd114: Instruction <= 32'h200834b8;
           10'd115: Instruction <= 32'hac0800d0;
           10'd116: Instruction <= 32'h20086be8;
           10'd117: Instruction <= 32'hac0800d4;
           10'd118: Instruction <= 32'h20084da4;
           10'd119: Instruction <= 32'hac0800d8;
           10'd120: Instruction <= 32'h20083aba;
           10'd121: Instruction <= 32'hac0800dc;
           10'd122: Instruction <= 32'h20080408;
           10'd123: Instruction <= 32'hac0800e0;
           10'd124: Instruction <= 32'h20086022;
           10'd125: Instruction <= 32'hac0800e4;
           10'd126: Instruction <= 32'h200826b7;
           10'd127: Instruction <= 32'hac0800e8;
           10'd128: Instruction <= 32'h2008797c;
           10'd129: Instruction <= 32'hac0800ec;
           10'd130: Instruction <= 32'h20082810;
           10'd131: Instruction <= 32'hac0800f0;
           10'd132: Instruction <= 32'h20081859;
           10'd133: Instruction <= 32'hac0800f4;
           10'd134: Instruction <= 32'h20084166;
           10'd135: Instruction <= 32'hac0800f8;
           10'd136: Instruction <= 32'h20084eb7;
           10'd137: Instruction <= 32'hac0800fc;
           10'd138: Instruction <= 32'h20086aca;
           10'd139: Instruction <= 32'hac080100;
           10'd140: Instruction <= 32'h2008722e;
           10'd141: Instruction <= 32'hac080104;
           10'd142: Instruction <= 32'h20081218;
           10'd143: Instruction <= 32'hac080108;
           10'd144: Instruction <= 32'h20087545;
           10'd145: Instruction <= 32'hac08010c;
           10'd146: Instruction <= 32'h20081373;
           10'd147: Instruction <= 32'hac080110;
           10'd148: Instruction <= 32'h2008707d;
           10'd149: Instruction <= 32'hac080114;
           10'd150: Instruction <= 32'h20084692;
           10'd151: Instruction <= 32'hac080118;
           10'd152: Instruction <= 32'h200800ea;
           10'd153: Instruction <= 32'hac08011c;
           10'd154: Instruction <= 32'h20084f8f;
           10'd155: Instruction <= 32'hac080120;
           10'd156: Instruction <= 32'h20081048;
           10'd157: Instruction <= 32'hac080124;
           10'd158: Instruction <= 32'h20081717;
           10'd159: Instruction <= 32'hac080128;
           10'd160: Instruction <= 32'h20087ae7;
           10'd161: Instruction <= 32'hac08012c;
           10'd162: Instruction <= 32'h20082d2d;
           10'd163: Instruction <= 32'hac080130;
           10'd164: Instruction <= 32'h200869f0;
           10'd165: Instruction <= 32'hac080134;
           10'd166: Instruction <= 32'h200832d4;
           10'd167: Instruction <= 32'hac080138;
           10'd168: Instruction <= 32'h20082ccb;
           10'd169: Instruction <= 32'hac08013c;
           10'd170: Instruction <= 32'h20080a6c;
           10'd171: Instruction <= 32'hac080140;
           10'd172: Instruction <= 32'h200872ab;
           10'd173: Instruction <= 32'hac080144;
           10'd174: Instruction <= 32'h20084b7c;
           10'd175: Instruction <= 32'hac080148;
           10'd176: Instruction <= 32'h20080d8d;
           10'd177: Instruction <= 32'hac08014c;
           10'd178: Instruction <= 32'h20081e3e;
           10'd179: Instruction <= 32'hac080150;
           10'd180: Instruction <= 32'h20087232;
           10'd181: Instruction <= 32'hac080154;
           10'd182: Instruction <= 32'h20080430;
           10'd183: Instruction <= 32'hac080158;
           10'd184: Instruction <= 32'h200804d8;
           10'd185: Instruction <= 32'hac08015c;
           10'd186: Instruction <= 32'h20087e6c;
           10'd187: Instruction <= 32'hac080160;
           10'd188: Instruction <= 32'h200800ba;
           10'd189: Instruction <= 32'hac080164;
           10'd190: Instruction <= 32'h200847a1;
           10'd191: Instruction <= 32'hac080168;
           10'd192: Instruction <= 32'h200878a6;
           10'd193: Instruction <= 32'hac08016c;
           10'd194: Instruction <= 32'h200846da;
           10'd195: Instruction <= 32'hac080170;
           10'd196: Instruction <= 32'h20082126;
           10'd197: Instruction <= 32'hac080174;
           10'd198: Instruction <= 32'h20084978;
           10'd199: Instruction <= 32'hac080178;
           10'd200: Instruction <= 32'h20085910;
           10'd201: Instruction <= 32'hac08017c;
           10'd202: Instruction <= 32'h2008460d;
           10'd203: Instruction <= 32'hac080180;
           10'd204: Instruction <= 32'h20084b7b;
           10'd205: Instruction <= 32'hac080184;
           10'd206: Instruction <= 32'h200836f6;
           10'd207: Instruction <= 32'hac080188;
           10'd208: Instruction <= 32'h20081e64;
           10'd209: Instruction <= 32'hac08018c;
           10'd210: Instruction <= 32'h200852ea;
           10'd211: Instruction <= 32'hac080190;
           10'd212: Instruction <= 32'h20087b94;
           10'd213: Instruction <= 32'hac080194;
           10'd214: Instruction <= 32'h20085ad7;
           10'd215: Instruction <= 32'hac080198;
           10'd216: Instruction <= 32'h20086d79;
           10'd217: Instruction <= 32'hac08019c;
           10'd218: Instruction <= 32'h20082fc0;
           10'd219: Instruction <= 32'hac0801a0;
           10'd220: Instruction <= 32'h20081817;
           10'd221: Instruction <= 32'hac0801a4;
           10'd222: Instruction <= 32'h2008387d;
           10'd223: Instruction <= 32'hac0801a8;
           10'd224: Instruction <= 32'h2008563f;
           10'd225: Instruction <= 32'hac0801ac;
           10'd226: Instruction <= 32'h20081e89;
           10'd227: Instruction <= 32'hac0801b0;
           10'd228: Instruction <= 32'h200845a7;
           10'd229: Instruction <= 32'hac0801b4;
           10'd230: Instruction <= 32'h2008624a;
           10'd231: Instruction <= 32'hac0801b8;
           10'd232: Instruction <= 32'h2008609a;
           10'd233: Instruction <= 32'hac0801bc;
           10'd234: Instruction <= 32'h20080a6d;
           10'd235: Instruction <= 32'hac0801c0;
           10'd236: Instruction <= 32'h20087a5b;
           10'd237: Instruction <= 32'hac0801c4;
           10'd238: Instruction <= 32'h20080f4e;
           10'd239: Instruction <= 32'hac0801c8;
           10'd240: Instruction <= 32'h20085b71;
           10'd241: Instruction <= 32'hac0801cc;
           10'd242: Instruction <= 32'h20086a88;
           10'd243: Instruction <= 32'hac0801d0;
           10'd244: Instruction <= 32'h2008656f;
           10'd245: Instruction <= 32'hac0801d4;
           10'd246: Instruction <= 32'h20083422;
           10'd247: Instruction <= 32'hac0801d8;
           10'd248: Instruction <= 32'h20082202;
           10'd249: Instruction <= 32'hac0801dc;
           10'd250: Instruction <= 32'h200841ed;
           10'd251: Instruction <= 32'hac0801e0;
           10'd252: Instruction <= 32'h20087f3a;
           10'd253: Instruction <= 32'hac0801e4;
           10'd254: Instruction <= 32'h20082313;
           10'd255: Instruction <= 32'hac0801e8;
           10'd256: Instruction <= 32'h20084b78;
           10'd257: Instruction <= 32'hac0801ec;
           10'd258: Instruction <= 32'h200860eb;
           10'd259: Instruction <= 32'hac0801f0;
           10'd260: Instruction <= 32'h20085560;
           10'd261: Instruction <= 32'hac0801f4;
           10'd262: Instruction <= 32'h20087783;
           10'd263: Instruction <= 32'hac0801f8;
           10'd264: Instruction <= 32'h200878bf;
           10'd265: Instruction <= 32'hac0801fc;
           10'd266: Instruction <= 32'h3c094000;
           10'd267: Instruction <= 32'h21290014;
           10'd268: Instruction <= 32'h8d230000;
           10'd269: Instruction <= 32'h20100080;
           10'd270: Instruction <= 32'h201101fc;
           10'd271: Instruction <= 32'h22320004;
           10'd272: Instruction <= 32'h00004020;
           10'd273: Instruction <= 32'h0111602a;
           10'd274: Instruction <= 32'h1180000d;
           10'd275: Instruction <= 32'h21090004;
           10'd276: Instruction <= 32'h0132602a;
           10'd277: Instruction <= 32'h11800008;
           10'd278: Instruction <= 32'h8d0a0000;
           10'd279: Instruction <= 32'h8d2b0000;
           10'd280: Instruction <= 32'h014b602a;
           10'd281: Instruction <= 32'h15800002;
           10'd282: Instruction <= 32'had2a0000;
           10'd283: Instruction <= 32'had0b0000;
           10'd284: Instruction <= 32'h21290004;
           10'd285: Instruction <= 32'h08000114;
           10'd286: Instruction <= 32'h21080004;
           10'd287: Instruction <= 32'h08000111;
           10'd288: Instruction <= 32'h3c094000;
           10'd289: Instruction <= 32'h21290014;
           10'd290: Instruction <= 32'h8d220000;
           10'd291: Instruction <= 32'h00431022;
           10'd292: Instruction <= 32'h200800c0;
           10'd293: Instruction <= 32'h20090710;
           10'd294: Instruction <= 32'had280000;
           10'd295: Instruction <= 32'h200800f9;
           10'd296: Instruction <= 32'had280004;
           10'd297: Instruction <= 32'h200800a4;
           10'd298: Instruction <= 32'had280008;
           10'd299: Instruction <= 32'h200800b0;
           10'd300: Instruction <= 32'had28000c;
           10'd301: Instruction <= 32'h20080099;
           10'd302: Instruction <= 32'had280010;
           10'd303: Instruction <= 32'h20080092;
           10'd304: Instruction <= 32'had280014;
           10'd305: Instruction <= 32'h20080082;
           10'd306: Instruction <= 32'had280018;
           10'd307: Instruction <= 32'h200800f8;
           10'd308: Instruction <= 32'had28001c;
           10'd309: Instruction <= 32'h20080080;
           10'd310: Instruction <= 32'had280020;
           10'd311: Instruction <= 32'h20080090;
           10'd312: Instruction <= 32'had280024;
           10'd313: Instruction <= 32'h20080088;
           10'd314: Instruction <= 32'had280028;
           10'd315: Instruction <= 32'h20080083;
           10'd316: Instruction <= 32'had28002c;
           10'd317: Instruction <= 32'h200800c6;
           10'd318: Instruction <= 32'had280030;
           10'd319: Instruction <= 32'h200800a1;
           10'd320: Instruction <= 32'had280034;
           10'd321: Instruction <= 32'h20080086;
           10'd322: Instruction <= 32'had280038;
           10'd323: Instruction <= 32'h2008008e;
           10'd324: Instruction <= 32'had28003c;
           10'd325: Instruction <= 32'h20080000;
           10'd326: Instruction <= 32'h11120003;
           10'd327: Instruction <= 32'h8d040000;
           10'd328: Instruction <= 32'h21080004;
           10'd329: Instruction <= 32'h08000146;
           10'd330: Instruction <= 32'h3c08ffff;
           10'd331: Instruction <= 32'h00084403;
           10'd332: Instruction <= 32'h2108ff9c;
           10'd333: Instruction <= 32'h3c094000;
           10'd334: Instruction <= 32'had280000;
           10'd335: Instruction <= 32'h3c08ffff;
           10'd336: Instruction <= 32'h00084403;
           10'd337: Instruction <= 32'had280004;
           10'd338: Instruction <= 32'h20080003;
           10'd339: Instruction <= 32'h3c094000;
           10'd340: Instruction <= 32'h21290008;
           10'd341: Instruction <= 32'had280000;
           10'd342: Instruction <= 32'h201b0000;
           10'd343: Instruction <= 32'h1000ffff;
           10'd344: Instruction <= 32'h20080001;
           10'd345: Instruction <= 32'h3c094000;
           10'd346: Instruction <= 32'h21290008;
           10'd347: Instruction <= 32'had280000;
           10'd348: Instruction <= 32'h200a0000;
           10'd349: Instruction <= 32'h136a0006;
           10'd350: Instruction <= 32'h214a0001;
           10'd351: Instruction <= 32'h136a0008;
           10'd352: Instruction <= 32'h214a0001;
           10'd353: Instruction <= 32'h136a000a;
           10'd354: Instruction <= 32'h214a0001;
           10'd355: Instruction <= 32'h136a000c;
           10'd356: Instruction <= 32'h2008000e;
           10'd357: Instruction <= 32'h00084200;
           10'd358: Instruction <= 32'h200b000f;
           10'd359: Instruction <= 32'h08000175;
           10'd360: Instruction <= 32'h2008000d;
           10'd361: Instruction <= 32'h00084200;
           10'd362: Instruction <= 32'h200b00f0;
           10'd363: Instruction <= 32'h08000175;
           10'd364: Instruction <= 32'h2008000b;
           10'd365: Instruction <= 32'h00084200;
           10'd366: Instruction <= 32'h200b0f00;
           10'd367: Instruction <= 32'h08000175;
           10'd368: Instruction <= 32'h20080007;
           10'd369: Instruction <= 32'h00084200;
           10'd370: Instruction <= 32'h200b0f00;
           10'd371: Instruction <= 32'h000b5900;
           10'd372: Instruction <= 32'h08000175;
           10'd373: Instruction <= 32'h004b6024;
           10'd374: Instruction <= 32'h11400004;
           10'd375: Instruction <= 32'h000c6102;
           10'd376: Instruction <= 32'h20010001;
           10'd377: Instruction <= 32'h01415022;
           10'd378: Instruction <= 32'h08000176;
           10'd379: Instruction <= 32'h000c4880;
           10'd380: Instruction <= 32'h21290710;
           10'd381: Instruction <= 32'h8d2a0000;
           10'd382: Instruction <= 32'h010a4020;
           10'd383: Instruction <= 32'h3c094000;
           10'd384: Instruction <= 32'h21290010;
           10'd385: Instruction <= 32'had280000;
           10'd386: Instruction <= 32'h237b0001;
           10'd387: Instruction <= 32'h20080003;
           10'd388: Instruction <= 32'h3c094000;
           10'd389: Instruction <= 32'h21290008;
           10'd390: Instruction <= 32'had280000;
           10'd391: Instruction <= 32'h200a0004;
           10'd392: Instruction <= 32'h176a0001;
           10'd393: Instruction <= 32'h201b0000;
           10'd394: Instruction <= 32'h03400008;
           10'd395: Instruction <= 32'h1000ffff;
           10'd396: Instruction <= 32'h03400008;
                
		      default: Instruction <= 32'h00000000;
		  endcase
endmodule
